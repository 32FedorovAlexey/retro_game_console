localparam FLY =     {32'b00000000_00000000_00000000_00000000,     //0
                       32'b00000000_00000000_00000000_00000000,     //1 
                       32'b00000000_00000000_00000000_00000000,     //
                       32'b00000000_00000000_00000000_00000000,     // 
                       32'b00000000_00000000_00000000_00000000,     // 
                       32'b00000000_00000000_00000000_00000000,     // 
                       32'b00000000_00000000_00000000_00000000,     //
                       32'b00000000_00000000_00000000_00000000,
                       32'b00000000_00000000_00000000_00000000,
                       32'b00000000_00000000_00000000_00000000,
                       32'b00000000_00000000_00000000_00000000,
		                 32'b00000000_00000000_00000000_00000000,
		                 32'b00000000_00000001_10000000_00000000,
		                 32'b00000000_00001111_11111000_00000000,
                       32'b00000000_11111111_11111111_00000000,
                       32'b00000111_11111110_01111111_11000000,
                       32'b00011111_11111100_00111111_11111000,
                       32'b00111111_11111110_01111111_11111100,
                       32'b00111000_00011110_01111100_00011100,
                       32'b01110000_00001111_11110000_00001110,
                       32'b01100000_00000111_11100000_00000110,
                       32'b01000000_00000011_11000000_00000010,
                       32'b01000000_00000011_11000000_00000010,
                       32'b00000000_00000001_10000000_00000000,
                       32'b00000000_00000001_10000000_00000000,
                       32'b00000000_00000001_10000000_00000000,
                       32'b00000000_00000001_10000000_00000000,
                       32'b00000000_00000001_10000000_00000000,
                       32'b00000000_00000001_10000000_00000000,
                       32'b00000000_00000001_10000000_00000000,
                       32'b00000000_00000001_10000000_00000000,
                       32'b00000000_00000001_10000000_00000000
		                }; 

localparam PLANE0 =  { 32'b00000000_00000001_00000000_00000000,
						     32'b00000000_00000001_00000000_00000000,
						     32'b00000000_00000011_10000000_00000000,
						     32'b00000000_00000011_10000000_00000000,
						     32'b00000000_00000111_11000000_00000000,
						     32'b00000000_00001111_11100000_00000000,
						     32'b00000000_00011111_11110000_00000000,
						     32'b00000000_00110001_10001100_00000000,
						     32'b00000000_01100001_10000110_00000000,
						     32'b00000000_11000001_10000011_00000000,
						     32'b00000001_10000001_10000001_10000000,
						     32'b00000011_00000001_10000000_11000000,
						     32'b00000110_00000001_10000000_01100000,
						     32'b00001100_00000001_10000000_00110000,
						     32'b00011100_00000001_10000000_00111000,
						     32'b00111000_00000001_10000000_00011100,
						     32'b00111000_00000001_10000000_00011100,
						     32'b00111000_00000001_10000000_00011100,
						     32'b00111111_11111111_11111111_11111100,
						     32'b00111111_11111111_11111111_01111100,
						     32'b00000000_00000001_10000000_00000000,
						     32'b00000000_00000001_10000000_00000000,
						     32'b00000000_00000001_10000000_00000000,
						     32'b00000000_00000001_10000000_00000000,
						     32'b00000000_00000001_10000000_00000000,
						     32'b00000000_00000011_11000000_00000000,
						     32'b00000000_00000111_11100000_00000000,
						     32'b00000000_00001111_11110000_00000000,
						     32'b00000000_00011111_11111000_00000000,
						     32'b00000000_00111111_11111100_00000000,
						     32'b00000000_00000000_00000000_00000000,
						     32'b00000000_00000000_00000000_00000000
						  } ;
localparam PLANE1 = {  32'b00000000_00000001_10000000_00000000,
						     32'b00000000_00000001_10000000_00000000,
						     32'b00000000_00000001_10000000_00000000,
						     32'b00000000_00000001_10000000_00000000,
						     32'b00000000_00000011_11000000_00000000,
						     32'b00000000_00000011_11000000_00000000,
						     32'b00000000_00000111_11100000_00000000,
						     32'b00000000_00001111_11110000_00000000,
						     32'b00000000_00001111_11110000_00000000,
						     32'b00000000_00011111_11111000_00000000,
						     32'b00000000_00011111_11111000_00000000,
						     32'b00010000_00011111_11111000_00001000,
						     32'b00111000_00011111_11111000_00011100,
						     32'b00111000_00111111_11111100_00011100,
						     32'b01111100_01111111_11111110_00111110,
						     32'b01111111_11111111_11111111_11111110,
						     32'b01111111_11111111_11111111_11111110,
						     32'b01111111_11111111_11111111_11111110,
						     32'b00011111_11111111_11111111_11111000,
						     32'b00000000_00000111_11100000_00000000,
						     32'b00000000_00000111_11100000_00000000,
						     32'b00000000_00000111_11100000_00000000,
						     32'b00000000_00001111_11110000_00000000,
						     32'b00000000_00011111_11111000_00000000,
						     32'b00000000_00000000_00000000_00000000,
						     32'b00000000_00000000_00000000_00000000,
						     32'b00000000_00000000_00000000_00000000,
						     32'b00000000_00000000_00000000_00000000,
						     32'b00000000_00000000_00000000_00000000,
						     32'b00000000_00000000_00000000_00000000,
						     32'b00000000_00000000_00000000_00000000,
						     32'b00000000_00000000_00000000_00000000
						  } ;						  
localparam BULLET = {   8'b00010000,
						      8'b00010000,
                        8'b00111000,
						      8'b00111000,
						      8'b00111000,
						      8'b00111000,
						      8'b01111100,
						      8'b11111110,
						  };						  