//  пробные символы
`define LETTER_30    {16'b1111111111111111, 16'b1111111111111111,16'b1110000000000111,16'b1111000000001111,16'b1101100000011011,16'b1100110000110011, 16'b1100011001100011,16'b1100001111000011,16'b1100000110000011,16'b1100001101100011,16'b1100110000110011,16'b1101100000011011,16'b1111000000001111,16'b1110000000000111,16'b1111111111111111,16'b1111111111111111}
`define LETTER_31    {16'hFF,16'hff,16'hff,16'hff,16'hff,16'hff,16'hff,16'hff,16'hff,16'hff,16'hff,16'hff,16'hff,16'hff,16'hff,16'hff}

// символы ASCII  цифра в названии это десятичный номер кода в таблице ASCII 
`define LETTER_32    {16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0}
`define LETTER_33    {16'd0,16'd24,16'd24,16'd24,16'd24,16'd24,16'd24,16'd24,16'd24,16'd0,16'd24,16'd24,16'd0,16'd0,16'd0,16'd0}
`define LETTER_34    {16'd0,16'd216,16'd216,16'd216,16'd216,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0 }
`define LETTER_35    {16'd408,16'd408,16'd408,16'd1020,16'd1020,16'd408,16'd408,16'd1020,16'd1020,16'd408,16'd408,16'd408,16'd0,16'd0,16'd0,16'd0 }
`define LETTER_36    {16'd0,16'd192,16'd192,16'd992,16'd1008,16'd240,16'd496,16'd992,16'd960,16'd1008,16'd496,16'd192,16'd192,16'd0,16'd0,16'd0 }
`define LETTER_37    {16'd0,16'd6192,16'd7288,16'd3788,16'd1740,16'd7116,16'd16376,16'd26544,16'd26304,16'd26336,16'd15472,16'd6192,16'd0,16'd0,16'd0,16'd0 }
`define LETTER_38    {16'd480,16'd1008,16'd824,16'd920,16'd440,16'd240,16'd240,16'd1016,16'd920,16'd792,16'd2040,16'd2032,16'd0,16'd0,16'd0,16'd0}
`define LETTER_39    {16'd0,16'd24,16'd24,16'd24,16'd24,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0}
`define LETTER_40    {16'd0,16'd48,16'd48,16'd24,16'd24,16'd24,16'd24,16'd24,16'd24,16'd24,16'd24,16'd48,16'd48,16'd0,16'd0,16'd0 }
`define LETTER_41    {16'd0,16'd48,16'd48,16'd96,16'd96,16'd96,16'd96,16'd96,16'd96,16'd96,16'd96,16'd48,16'd48,16'd0,16'd0,16'd0 }
`define LETTER_42    {16'd48,16'd252,16'd252,16'd120,16'd252,16'd204,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0 }
`define LETTER_43    {16'd0,16'd0,16'd0,16'd0,16'd96,16'd96,16'd504,16'd504,16'd96,16'd96,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0 }
`define LETTER_44    {16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd24,16'd24,16'd16,16'd8,16'd0,16'd0}
`define LETTER_45    {16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd504,16'd504,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0}
`define LETTER_46    {16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd24,16'd24,16'd0,16'd0,16'd0,16'd0}
`define LETTER_47    {16'd192,16'd192,16'd224,16'd96,16'd112,16'd48,16'd48,16'd56,16'd24,16'd28,16'd12,16'd12,16'd0,16'd0,16'd0,16'd0}
`define LETTER_48    {16'd0,16'd496,16'd1016,16'd984,16'd984,16'd984,16'd856,16'd888,16'd888,16'd888,16'd1016,16'd496,16'd0,16'd0,16'd0,16'd0}
`define LETTER_49    {16'd0,16'd192,16'd224,16'd240,16'd240,16'd192,16'd192,16'd192,16'd192,16'd192,16'd1008,16'd1008,16'd0,16'd0,16'd0,16'd0}

`define LETTER_50    {16'd0,16'd240,16'd504,16'd408,16'd384,16'd384,16'd448,16'd224,16'd112,16'd120,16'd504,16'd504,16'd0,16'd0,16'd0,16'd0}
`define LETTER_51    {16'd0,16'd240,16'd504,16'd408,16'd384,16'd448,16'd192,16'd448,16'd384,16'd408,16'd504,16'd240,16'd0,16'd0,16'd0,16'd0}
`define LETTER_52    {16'd0,16'd384,16'd448,16'd480,16'd496,16'd440,16'd408,16'd1016,16'd1016,16'd384,16'd384,16'd384,16'd0,16'd0,16'd0,16'd0}
`define LETTER_53    {16'd0,16'd504,16'd504,16'd24,16'd24,16'd248,16'd504,16'd384,16'd384,16'd408,16'd504,16'd240,16'd0,16'd0,16'd0,16'd0}
`define LETTER_54    {16'd0,16'd240,16'd504,16'd408,16'd24,16'd248,16'd504,16'd408,16'd408,16'd408,16'd504,16'd240,16'd0,16'd0,16'd0,16'd0}
`define LETTER_55    {16'd0,16'd1016,16'd1016,16'd768,16'd896,16'd448,16'd224,16'd96,16'd96,16'd96,16'd96,16'd96,16'd0,16'd0,16'd0,16'd0}
`define LETTER_56    {16'd0,16'd240,16'd504,16'd408,16'd408,16'd240,16'd504,16'd408,16'd408,16'd408,16'd504,16'd240,16'd0,16'd0,16'd0,16'd0}
`define LETTER_57    {16'd0,16'd240,16'd504,16'd408,16'd408,16'd504,16'd496,16'd384,16'd384,16'd408,16'd504,16'd240,16'd0,16'd0,16'd0,16'd0}
`define LETTER_58    {16'd0,16'd0,16'd0,16'd0,16'd24,16'd24,16'd0,16'd0,16'd0,16'd0,16'd24,16'd24,16'd0,16'd0,16'd0,16'd0}
`define LETTER_59    {16'd0,16'd0,16'd0,16'd0,16'd24,16'd24,16'd0,16'd0,16'd0,16'd0,16'd24,16'd24,16'd16,16'd8,16'd0,16'd0}

`define LETTER_60    {16'd0,16'd0,16'd0,16'd3840,16'd4032,16'd1008,16'd124,16'd124,16'd1008,16'd4032,16'd3840,16'd0,16'd0,16'd0,16'd0,16'd0}
`define LETTER_61    {16'd0,16'd0,16'd0,16'd0,16'd504,16'd504,16'd0,16'd0,16'd504,16'd504,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0}
`define LETTER_62    {16'd0,16'd0,16'd0,16'd60,16'd252,16'd1008,16'd3968,16'd3968,16'd1008,16'd252,16'd60,16'd0,16'd0,16'd0,16'd0,16'd0}
`define LETTER_63    {16'd0,16'd240,16'd504,16'd408,16'd384,16'd448,16'd224,16'd96,16'd96,16'd0,16'd96,16'd96,16'd0,16'd0,16'd0,16'd0}
`define LETTER_64    {16'd0,16'd8160,16'd16368,16'd28728,16'd26520,16'd28632,16'd27864,16'd27864,16'd27864,16'd27864,16'd32728,16'd16280,16'd56,16'd16368,16'd16352,16'd0}
`define LETTER_65    {16'd0,16'd480,16'd1008,16'd1848,16'd1560,16'd1560,16'd2040,16'd2040,16'd1560,16'd1560,16'd1560,16'd1560,16'd0,16'd0,16'd0,16'd0}
`define LETTER_66    {16'd0,16'd1016,16'd2040,16'd1560,16'd1560,16'd2040,16'd1016,16'd1560,16'd1560,16'd1560,16'd2040,16'd1016,16'd0,16'd0,16'd0,16'd0}
`define LETTER_67    {16'd0,16'd992,16'd2032,16'd1584,16'd48,16'd48,16'd48,16'd48,16'd48,16'd1584,16'd2032,16'd992,16'd0,16'd0,16'd0,16'd0}
`define LETTER_68    {16'd0,16'd2032,16'd4080,16'd3120,16'd3120,16'd3120,16'd3120,16'd3120,16'd3120,16'd3120,16'd4080,16'd2032,16'd0,16'd0,16'd0,16'd0}
`define LETTER_69    {16'd0,16'd1008,16'd1008,16'd48,16'd48,16'd1008,16'd1008,16'd48,16'd48,16'd48,16'd1008,16'd1008,16'd0,16'd0,16'd0,16'd0}

`define LETTER_70    {16'd0,16'd1008,16'd1008,16'd48,16'd48,16'd1008,16'd1008,16'd48,16'd48,16'd48,16'd48,16'd48,16'd0,16'd0,16'd0,16'd0}
`define LETTER_71    {16'd0,16'd992,16'd2032,16'd1584,16'd48,16'd48,16'd1840,16'd1840,16'd1584,16'd1584,16'd2032,16'd992,16'd0,16'd0,16'd0,16'd0}
`define LETTER_72    {16'd0,16'd1560,16'd1560,16'd1560,16'd1560,16'd2040,16'd2040,16'd1560,16'd1560,16'd1560,16'd1560,16'd1560,16'd0,16'd0,16'd0,16'd0}
`define LETTER_73    {16'd0, 16'd120, 16'd120, 16'd48, 16'd48, 16'd48, 16'd48, 16'd48, 16'd48, 16'd48, 16'd120, 16'd120, 16'd0,16'd0,16'd0,16'd0}
`define LETTER_74    {16'd0,16'd480,16'd480,16'd192,16'd192,16'd192,16'd192,16'd192,16'd192,16'd204,16'd252,16'd120,16'd0,16'd0,16'd0,16'd0}
`define LETTER_75    {16'd0,16'd1560,16'd1816,16'd920,16'd472,16'd248,16'd120,16'd248,16'd472,16'd920,16'd1816,16'd1560,16'd0,16'd0,16'd0,16'd0}
`define LETTER_76    {16'd0,16'd24,16'd24,16'd24,16'd24,16'd24,16'd24,16'd24,16'd24,16'd24,16'd504,16'd04,16'd0,16'd0,16'd0,16'd0}
`define LETTER_77    {16'd0,16'd6168,16'd7224,16'd7800,16'd8184,16'd7128,16'd6552,16'd6168,16'd6168,16'd6168,16'd6168,16'd6168,16'd0,16'd0,16'd0,16'd0}
`define LETTER_78    {16'd0,16'd3096,16'd3128,16'd3192,16'd3320,16'd3576,16'd3544,16'd4056,16'd3992,16'd3864,16'd3608,16'd3096,16'd0,16'd0,16'd0,16'd0}
`define LETTER_79    {16'd0,16'd2016,16'd4080,16'd3120,16'd3120,16'd3120,16'd3120,16'd3120,16'd3120,16'd3120,16'd4080,16'd2016,16'd0,16'd0,16'd0,16'd0}

`define LETTER_80    {16'd0,16'd504,16'd1016,16'd792,16'd792,16'd792,16'd1016,16'd504,16'd24,16'd24,16'd24,16'd24,16'd0,16'd0,16'd0,16'd0}
`define LETTER_81    {16'd0,16'd2016,16'd4080,16'd3120,16'd3120,16'd3120,16'd3120,16'd3120,16'd3120,16'd3632,16'd4080,16'd8160,16'd0,16'd0,16'd0,16'd0}
`define LETTER_82    {16'd0,16'd1016,16'd2040,16'd1560,16'd1560,16'd2040,16'd1016,16'd1560,16'd1560,16'd1560,16'd1560,16'd1560,16'd0,16'd0,16'd0,16'd0}
`define LETTER_83    {16'd0,16'd1008,16'd2040,16'd1560,16'd24,16'd1016,16'd2032,16'd1536,16'd1536,16'd1560,16'd2040,16'd1008,16'd0,16'd0,16'd0,16'd0}
`define LETTER_84    {16'd0,16'd2040,16'd2040,16'd192,16'd192,16'd192,16'd192,16'd192,16'd192,16'd192,16'd192,16'd192,16'd0,16'd0,16'd0,16'd0}
`define LETTER_85    {16'd0,16'd3120,16'd3120,16'd3120,16'd3120,16'd3120,16'd3120,16'd3120,16'd3120,16'd3120,16'd4080,16'd2016,16'd0,16'd0,16'd0,16'd0}
`define LETTER_86    {16'd0,16'd3120,16'd3120,16'd3120,16'd3120,16'd3120,16'd3120,16'd3120,16'd3696,16'd2016,16'd960,16'd384,16'd0,16'd0,16'd0,16'd0}
`define LETTER_87    {16'd0,16'd6168,16'd6168,16'd6168,16'd6552,16'd6552,16'd6552,16'd6552,16'd6552,16'd8184,16'd4080,16'd1632,16'd0,16'd0,16'd0,16'd0}
`define LETTER_88    {16'd0,16'd1560,16'd1848,16'd816,16'd1008,16'd480,16'd192,16'd480,16'd1008,16'd816,16'd1848,16'd1560,16'd0,16'd0,16'd0,16'd0}
`define LETTER_89    {16'd0,16'd1560,16'd1848,16'd816,16'd1008,16'd480,16'd192,16'd192,16'd192,16'd192,16'd192,16'd192,16'd0,16'd0,16'd0,16'd0}

`define LETTER_90    {16'd0,16'd4092,16'd4092,16'd1792,16'd896,16'd448,16'd192,16'd224,16'd112,16'd56,16'd4092,16'd4092,16'd0,16'd0,16'd0,16'd0}

/*
localparam logic [0:60][15:0][15:0] bitmap = {   `LETTER_32,`LETTER_33,`LETTER_32,`LETTER_33,`LETTER_34,`LETTER_35,`LETTER_36,`LETTER_37,`LETTER_38,`LETTER_39,  
                                                 `LETTER_40,`LETTER_41,`LETTER_42,`LETTER_43,`LETTER_44,`LETTER_45,`LETTER_46,`LETTER_47,`LETTER_48,`LETTER_49,     
                                                 `LETTER_50,`LETTER_51,`LETTER_52,`LETTER_53,`LETTER_54,`LETTER_55,`LETTER_56,`LETTER_57,`LETTER_58,`LETTER_59,     
                                                 `LETTER_60,`LETTER_61,`LETTER_62,`LETTER_63,`LETTER_64,`LETTER_65,`LETTER_66,`LETTER_67,`LETTER_68,`LETTER_69,     
                                                 `LETTER_70,`LETTER_71,`LETTER_72,`LETTER_73,`LETTER_74,`LETTER_75,`LETTER_76,`LETTER_77,`LETTER_78,`LETTER_79,
                                                 `LETTER_80,`LETTER_81,`LETTER_82,`LETTER_83,`LETTER_84,`LETTER_85,`LETTER_86,`LETTER_87,`LETTER_88,`LETTER_89,
                                                 `LETTER_90}; 

localparam logic [0:9][15:0][15:0] bitmap_n = {   `LETTER_48,`LETTER_49,`LETTER_50,`LETTER_51,`LETTER_52,`LETTER_53,`LETTER_54,`LETTER_55,`LETTER_56,`LETTER_57}; 
*/       