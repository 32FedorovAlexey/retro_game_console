
module retro_game  ( 
                    input  clk,
						  input  key_right,
						  input  key_left,
						  input  key_fire,
						  output v_sync,
						  output h_sync,
						  output r_pin,
						  output g_pin,
						  output b_pin
						 );
						 
						 
         vga  vga_i
                   ( 
						  .clk(clk),
                    .rst(1'b0),                            // сигнал нужен для моделирования при имплементации можно установить в "0" 
                    .h_sync(h_sync),
                    .v_sync(v_sync),
                    .x(x),
                    .y(y)
          );						 
						 
    wire [9:0] x,y;
	 reg        r,g,b;
	 reg  [7:0] count_1, count_2;
	 
	 
	 
	 
	  
	 // задаем частоту просчета сцены 
	 
	 logic tik;
	 
    low_clock  #(.F_CLK_SLOW(20))
	      low_clock_i 
                   (
						  .clk(clk),
                    .rst(1'b0),
                    .clk_slow(),
                    .one_pulse(tik)
                    );

// триггер попаданий
	 reg        was_hit;  
	 wire  crash = flyer_g & bullet_r ;
	
   always_ff @(posedge clk) 
	  if (tik) was_hit <= 1'b0;
	  else if (crash) was_hit <= 1'b1;
 	
	// главный цикл геймплея
	  
	 always_ff @(posedge clk)
	 if(tik)
	   begin
		// движение коробля пришельцнв 
         f_x_pos   <= (f_dir_mov)?  f_x_pos - 5 : f_x_pos + 5;
	      if (f_x_pos < 10'd6)   f_dir_mov <= 1'b0;	
	      if (f_x_pos > 10'd600) f_dir_mov <= 1'b1;	
      	
	
   	// движение самолета  
        if (( ~key_left ) & ( p_x_pos > 11'd1))   p_x_pos <= p_x_pos - 2;
		  if (( ~key_right) & ( p_x_pos < 11'd608)) p_x_pos <= p_x_pos + 2;

	   	// движение снаряда
	     if (~key_fire & ~bullet_mov) begin                // нажали кнопку fire
		    bullet_mov <=1'b1;	
          count_1 <= count_1 + 1;	
	       if (count_1[3:0] == 4'h9)
			    count_1<= count_1 + 4'h7;		                // двоично-десятичная корекция 
			end
		   //else 
			
			if (was_hit & bullet_mov) begin                  //снаряд встретился с кораблем пришельцев 
			   count_2 <= count_2 + 1;
				if (count_2[3:0] == 4'h9)
			     count_2<= count_2 + 4'h7;	                // двоично-десятичная корекция 
			end 			  
			
		  if ((bullet_y < 20) | was_hit) begin               // вышли за пределы экрана или встретились с кораблем пришельцев
		    bullet_mov <= 1'b0;
  		//	 bullet_y <= p_y_pos ;                            // возвращаем  снаряд на корабль
		//	 bullet_x <= p_x_pos + 13;
		  end

		  if (bullet_mov) 
		    bullet_y <= bullet_y - 5;                       // движение снаряда
		  else begin  
		  	 bullet_y <= p_y_pos ;                           // возвращаем  снаряд на корабль
			 bullet_x <= p_x_pos + 12;
		  end
	  
	   end 	 

		
     // wire r_sqr = ((x > 13) & (x < 18) & (y > 80) & (y < 130)) ? 1'b1 : 1'b0 ; // красный квадрат
	  
	// счетчик выстрелов 
 logic shot_r,shot_g, shot_b;
    numbers  shot	 
           ( .x(x),
             .y(y),
				 .data({count_1[3:0],count_1[7:4]}),                               //  выводимые цифры  
             .pos_x(10'd600),
             .pos_y(10'd30),
             .collor(3'b011),
             
             .r(shot_r), 
             .g(shot_g), 
             .b(shot_b)
            );	
	 
	 // надпись "SHOT"
	 	logic text1_r,text1_g,text1_b;
    
	 text #(.L(5), 
         .data({8'd53, 8'd42, 8'd49, 8'd54, 8'd28 })
        )
            text_shot (
                    .x(x),
				        .y(y),
				        .pos_x(10'd520),  
						  .pos_y(10'd30),
						  .collor(3'b011),
						  .r(text1_r),
                    .g(text1_g),
						  .b(text1_b)

						  );			
 

	 
	 // счетчик попаданий
	 logic hit_r,hit_g,hit_b;
    numbers  hit	 
           ( .x(x),
             .y(y),
				 .data({count_2[3:0],count_2[7:4]}),                               // выводимые цифры  
             .pos_x(10'd600),
             .pos_y(10'd46),
             .collor(3'b100),
             
             .r(hit_r), 
             .g(hit_g), 
             .b(hit_b)
            );				
	
	
 
	 // надпись "HIT"
	 logic text2_r,text2_g,text2_b;	
     text #(.L(4), 
         .data({8'd42, 8'd43, 8'd54, 8'd28 })
        )
            text_hit (
                    .x(x),
				        .y(y),
				        .pos_x(10'd536),  
						  .pos_y(10'd46),
						  .collor(3'b100),
						  .r(text2_r),
                    .g(text2_g),
						  .b(text2_b)
						  );			

	 
	 logic       plane_r,plane_g,plane_b;
	 logic [9:0] p_x_pos = 10'd320;
	 logic [9:0] p_y_pos = 10'd440;
	       

    sprite  #(.SIZE(32), 
	           .MASK(
				       {32'b00000000_00000001_00000000_00000000,
						  32'b00000000_00000001_00000000_00000000,
						  32'b00000000_00000011_10000000_00000000,
						  32'b00000000_00000011_10000000_00000000,
						  32'b00000000_00000111_11000000_00000000,
						  32'b00000000_00001111_11100000_00000000,
						  32'b00000000_00011111_11110000_00000000,
						  32'b00000000_00110001_10001100_00000000,
						  32'b00000000_01100001_10000110_00000000,
						  32'b00000000_11000001_10000011_00000000,
						  32'b00000001_10000001_10000001_10000000,
						  32'b00000011_00000001_10000000_11000000,
						  32'b00000110_00000001_10000000_01100000,
						  32'b00001100_00000001_10000000_00110000,
						  32'b00011100_00000001_10000000_00111000,
						  32'b00111000_00000001_10000000_00011100,
						  32'b00111000_00000001_10000000_00011100,
						  32'b00111000_00000001_10000000_00011100,
						  32'b00111111_11111111_11111111_11111100,
						  32'b00111111_11111111_11111111_01111100,
						  32'b00000000_00000001_10000000_00000000,
						  32'b00000000_00000001_10000000_00000000,
						  32'b00000000_00000001_10000000_00000000,
						  32'b00000000_00000001_10000000_00000000,
						  32'b00000000_00000001_10000000_00000000,
						  32'b00000000_00000011_11000000_00000000,
						  32'b00000000_00000111_11100000_00000000,
						  32'b00000000_00001111_11110000_00000000,
						  32'b00000000_00011111_11111000_00000000,
						  32'b00000000_00111111_11111100_00000000,
						  32'b00000000_00000000_00000000_00000000,
						  32'b00000000_00000000_00000000_00000000
						  }))
						  
	           plane(
	                 .x(x),
				        .y(y),
				        .pos_x(p_x_pos),
						  .pos_y(p_y_pos),
						  .collor(3'b100),
						  .r(plane_r),
                    .g(plane_g),
						  .b(plane_b)
						 );	
						 
			logic [9:0] bullet_x, bullet_y;
			logic       bullet_mov, bullet_r,bullet_g,bullet_b;
			
	sprite  #(.SIZE(8), 
	           .MASK(
				       { 8'b00010000,
						   8'b00010000,
                     8'b00111000,
						   8'b00111000,
						   8'b00111000,
						   8'b00111000,
						   8'b01111100,
						   8'b11111110,
						  }))
						  
	           bullet(
	                 .x(x),
				        .y(y),
				        .pos_x(bullet_x),
						  .pos_y(bullet_y),
						  .collor(3'b100),
						  .r(bullet_r),
                    .g(bullet_g),
						  .b(bullet_b)
						 );	
						 					 
						 
				logic       flyer_r,flyer_g,flyer_b;
	         logic [9:0] f_x_pos;                                 // координата х корабля пришельцев
            logic       f_dir_mov;                               // Нарпавление движения 0 в право 1 в лево     
   			
				sprite  #(.SIZE(32), 
	           .MASK(
				       {32'b00000000_00000000_00000000_00000000,     //0
						  32'b00000000_00000000_00000000_00000000,     //1 
						  32'b00000000_00000000_00000000_00000000,     //
						  32'b00000000_00000000_00000000_00000000,     // 
						  32'b00000000_00000000_00000000_00000000,     // 
						  32'b00000000_00000000_00000000_00000000,     // 
						  32'b00000000_00000000_00000000_00000000,     //
						  32'b00000000_00000000_00000000_00000000,
						  32'b00000000_00000000_00000000_00000000,
						  32'b00000000_00000000_00000000_00000000,
						  32'b00000000_00000000_00000000_00000000,
						  32'b00000000_00000000_00000000_00000000,
						  32'b00000000_00000001_10000000_00000000,
						  32'b00000000_00001111_11111000_00000000,
						  32'b00000000_11111111_11111111_00000000,
						  32'b00000111_11111110_01111111_11000000,
						  32'b00011111_11111100_00111111_11111000,
						  32'b00111111_11111110_01111111_11111100,
						  32'b00111000_00011110_01111100_00011100,
						  32'b01110000_00001111_11110000_00001110,
						  32'b01100000_00000111_11100000_00000110,
						  32'b01000000_00000011_11000000_00000010,
						  32'b01000000_00000011_11000000_00000010,
						  32'b00000000_00000001_10000000_00000000,
						  32'b00000000_00000001_10000000_00000000,
						  32'b00000000_00000001_10000000_00000000,
						  32'b00000000_00000001_10000000_00000000,
						  32'b00000000_00000001_10000000_00000000,
						  32'b00000000_00000001_10000000_00000000,
						  32'b00000000_00000001_10000000_00000000,
						  32'b00000000_00000001_10000000_00000000,
						  32'b00000000_00000001_10000000_00000000
						  }))
						  
	           flyer(
	                 .x(x),
				        .y(y),
				        .pos_x(f_x_pos),
						  .pos_y(80),
						  .collor(3'b010),
						  .r(flyer_r),
                    .g(flyer_g),
						  .b(flyer_b)
						 );	
 						 
/*	logic text_r, text_g, text_b;
	
  text #(.L(14), 
         .data({8'd35, 8'd46, 8'd39, 8'd58, 8'd39, 8'd59, 8'd2, 8'd40, 8'd39, 8'd38, 8'd49, 8'd52, 8'd49, 8'd56})
        )
            text_1 (
                    .x(x),
				        .y(y),
				        .pos_x(250), //250
						  .pos_y(50),
						  .collor(3'b111),
						  .r(text_r),
                    .g(text_g),
						  .b(text_b)

						  );			
*/

	logic lw1;					  
	/*line line_1(
	            .clk(clk),
					.x(x),
					.y(y),
					.x1(10'd280),
					.x2(10'd320),
					.y1(10'd150),
					.y2(10'd150),
					.white(lw1)
					);					  
*/
		logic lw2;					  
	/*line line_2(
	            .clk(clk),
					.x(x),
					.y(y),
					.x1(10'd280),
					.x2(10'd350),
					.y1(10'd150),
					.y2(10'd200),
					.white(lw2)
					);					 
	*/
	logic lw3;					  
	/*line line_3(
	            .clk(clk),
					.x(x),
					.y(y),
					.x1(10'd320),
					.x2(10'd350),
					.y1(10'd150),
					.y2(10'd200),
					.white(lw3)
					);					  
  		*/		
  			
   assign r_pin = plane_r | flyer_r | bullet_r | shot_r | hit_r  | text1_r | text2_r | lw1 | lw2 | lw3 ; 
   assign g_pin = plane_g | flyer_g | bullet_g | shot_g | hit_g  | text1_g | text2_g | lw1 | lw2 | lw3 ; 
   assign b_pin = plane_b | flyer_b | bullet_b | shot_b | hit_b  | text1_b | text2_b | lw1 | lw2 | lw3 ; 
  
  
  
endmodule 
						 